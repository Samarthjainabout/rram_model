* ReRAM Step Pulse Time Analysis

* Default values
.param VSTEP=1.8
.param PW=100n

V1 TE 0 PULSE(0 {VSTEP} 0 1n 1n {PW} {2*PW})

XR0 TE 0 sky130_fd_pr_reram__reram_cell Tfilament_0=3.8e-9

.tran 0.1n 2u

.include /content/rram_model/ngspice/sky130_fd_pr_reram__reram_cell.spice

.control
set filetype=ascii

alter .param PW=10n
run
write pw_10n.raw

alter .param PW=50n
run
write pw_50n.raw

alter .param PW=100n
run
write pw_100n.raw

alter .param PW=500n
run
write pw_500n.raw

alter .param PW=1u
run
write pw_1u.raw

.endc

.end
