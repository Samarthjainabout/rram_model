ReRAM Example

.param VSTEP=1.8
.param PW=100n

V1 TE 0 PULSE(0 {VSTEP} 0 1n 1n {PW} {2*PW})

XR0 TE 0 sky130_fd_pr_reram__reram_cell Tfilament_0=3.8e-9

.tran 0.1n 2u
.step param PW list 10n 50n 100n 500n 1u

.inc /foss/pdks/sky130B/libs.tech/ngspice/sky130_fd_pr_reram__reram_cell.spice

.control
set filetype=ascii
.endc

.end
